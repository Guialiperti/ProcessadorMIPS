library ieee;
use ieee.std_logic_1164.all;

entity muxGenerico2_1bit is
    generic (
        -- Total de bits das entradas e saidas
        larguraDados    : natural  :=   8
    );
    port (
        entradaA    : in  std_logic;
        entradaB    : in  std_logic;
        seletor     : in  std_logic;
        saida       : out std_logic
    );
end entity;

architecture comportamento of muxGenerico2_1bit is
begin
  -- Para sintetizar lógica combinacional usando um processo,
  --  todas as entradas do modulo devem aparecer na lista de sensibilidade.
    process(entradaA, entradaB, seletor) is
    begin
        if(seletor='0') then
            saida <= entradaA;
        else
            saida <= entradaB;
        end if;
    end process;
end architecture;